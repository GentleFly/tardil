
(* dont_touch="true" *)
module inv (
  input i,
  output o
);
  assign o = ~i;
endmodule

